** sch_path: /home/uri/p/tt10-simon-game/xschem/ring_osc.sch
**.subckt ring_osc
V1 VSS 0 0
V2 VDD VSS 3.3
x1 net13 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x2 net2 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x3 net3 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x4 net4 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x5 net5 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x6 net6 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x7 net1 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x8 net7 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x9 net8 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x10 net9 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x11 net10 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x12 net11 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x13 net12 clk_out VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x14 en clk_out net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
x15 VDD en VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
C1 net13 VSS 2f m=1
C2 net2 VSS 2f m=1
C3 net3 VSS 2f m=1
C4 net4 VSS 2f m=1
C5 net5 VSS 2f m=1
C6 net6 VSS 2f m=1
C7 net1 VSS 2f m=1
C8 net7 VSS 2f m=1
C9 net8 VSS 2f m=1
C10 net9 VSS 2f m=1
C11 net10 VSS 2f m=1
C12 net11 VSS 2f m=1
C13 net12 VSS 2f m=1
**** begin user architecture code

.include design.ngspice
.lib sm141064.ngspice typical
.include gf180mcu_fd_sc_mcu7t5v0.spice

.control
save all
tran 10p 100n
write ring_osc.raw
meas tran tdiff TRIG clk_out VAL=3 RISE=20 TARG clk_out VAL=3 RISE=21
let freq_mhz = (1 / (tdiff) / 1e6)
print freq_mhz
plot clk_out
.endc


**** end user architecture code
**.ends
.end
